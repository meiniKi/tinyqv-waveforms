`default_nettype none
`timescale 1ns / 1ps

/* This testbench just instantiates the module and makes some convenient wires
   that can be driven / tested by the cocotb test.py.
*/
module tb ();

  // Dump the signals to a VCD file. You can view it with gtkwave or surfer.
  initial begin
    $dumpfile("tb.vcd");
    $dumpvars(0, tb);
    #1;
  end

  // Wire up the inputs and outputs:
  reg clk;
  reg rst_n;
  reg ena;
  reg [7:0] ui_in;
  reg [7:0] uio_in;
  wire [7:0] uo_out;
  wire [7:0] uio_out;
  wire [7:0] uio_oe;
`ifdef GL_TEST
  wire VPWR = 1'b1;
  wire VGND = 1'b0;
`endif

  tt_um_tqv_peripheral_harness test_harness (

      // Include power ports for the Gate Level test:
`ifdef GL_TEST
      .VPWR(VPWR),
      .VGND(VGND),
`endif

      .ui_in  (ui_in),    // Dedicated inputs
      .uo_out (uo_out),   // Dedicated outputs
      .uio_in (uio_in),   // IOs: Input path
      .uio_out(uio_out),  // IOs: Output path
      .uio_oe (uio_oe),   // IOs: Enable path (active high: 0=input, 1=output)
      .ena    (ena),      // enable - goes high when design is selected
      .clk    (clk),      // clock
      .rst_n  (rst_n)     // not reset
  );

  (* keep *) wire tst_cs;
  (* keep *) wire tst_sd;
  (* keep *) wire tst_sck;
  (* keep *) wire tst_dc;

  assign tst_cs   = uo_out[3];
  assign tst_sd   = uo_out[2];
  assign tst_sck  = uo_out[1];
  assign tst_dc   = uo_out[4];

`ifdef MODEL
  ssd1306_spi4 i_ssd1306_spi4 (
    .cs_in  ( uo_out[3] ),
    .sdi_i  ( uo_out[2] ),
    .sck_i  ( uo_out[1] ),
    .dc_i   ( uo_out[4] )
  );
`endif



endmodule
